library verilog;
use verilog.vl_types.all;
entity Maquina_de_refri_vlg_vec_tst is
end Maquina_de_refri_vlg_vec_tst;
